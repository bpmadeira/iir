https://github.com/oscimp/oscimpDigital
